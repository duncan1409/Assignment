module mx2_32bits(

);
endmodule