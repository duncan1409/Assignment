module ha(
	input a, b,
	output y
	);
	
	_and2 ad20 (
		.a(a),
		b.(b),
		y.(y)
	
endmodule