module cla4_ov(

);
endmodule