`timescale 1ns/100ps
module tb_alu4 (

);
endmodule