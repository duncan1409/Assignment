module cal_flags4(

);
endmodule