module mx8_32bits(

);
endmodule