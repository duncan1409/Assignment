module ha (
	input a, b,
	output co, s
	);
	
	_and2 ad20 (
		.a(a),
		.b(b),
		.y(co)
		);
	
	_or2 or20 (
		.a(a),
		.b(b),
		.y(s)
		);
	
endmodule
