module mx2_4bits(

);
endmodule