module (clk, reset_n, Ta, Tal, Tb, Tbl, La, Lb)
  input clk, reset_n, Ta, Tal, Tb, Tbl;
  output [1:0] La, Lb;

endmodule