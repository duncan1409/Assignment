module (clk, reset_n, Ta, Tb, La, Lb);
  input clk, reset_n, Ta, Tb;
  output La, Lb;

endmodule