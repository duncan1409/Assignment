module cla32_ov(

);
endmodule