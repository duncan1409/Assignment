module mx8_4bits(

);
endmodule