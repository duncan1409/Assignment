module cal_flags32(

);
endmodule