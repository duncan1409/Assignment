module alu32(

);
endmodule