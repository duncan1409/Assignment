module alu4 (

);
endmodule